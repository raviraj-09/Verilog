module Half_Substractor(input A, B, output Dif, bow);
assign dif = A^B;
assign bow = ~A&B;
endmodule
